* SPICE3 file created from INVX1_new.ext - technology: scmos

.subckt INVX1_new A Y vdd gnd
M1000 Y gnd vdd vdd pfet w=2.1u l=0.6u
+  ad=3.15p pd=7.2u as=3.15p ps=7.2u
M1001 Y A gnd Gnd nfet w=3.9u l=0.6u
+  ad=5.85p pd=10.8u as=5.85p ps=10.8u
C0 gnd vdd 2.89fF
C1 gnd Gnd 4.57fF
C2 vdd Gnd 6.00fF
.ends

X100 A Z VDD GND INVX1_new
.end