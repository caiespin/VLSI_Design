magic
tech scmos
timestamp 1551173462
<< nwell >>
rect 170 -4 194 25
<< ntransistor >>
rect 181 -17 183 -13
<< ptransistor >>
rect 181 2 183 14
<< ndiffusion >>
rect 180 -17 181 -13
rect 183 -17 184 -13
<< pdiffusion >>
rect 180 2 181 14
rect 183 2 184 14
<< ndcontact >>
rect 176 -17 180 -13
rect 184 -17 188 -13
<< pdcontact >>
rect 176 2 180 14
rect 184 2 188 14
<< psubstratepcontact >>
rect 176 -46 180 -42
<< nsubstratencontact >>
rect 176 18 180 22
<< polysilicon >>
rect 181 14 183 16
rect 181 -13 183 2
rect 181 -19 183 -17
<< polycontact >>
rect 177 -8 181 -4
<< metal1 >>
rect 169 23 194 27
rect 176 22 180 23
rect 176 14 180 18
rect 184 -4 188 2
rect 168 -8 177 -4
rect 184 -8 196 -4
rect 184 -13 188 -8
rect 176 -42 180 -17
rect 169 -50 194 -46
<< labels >>
rlabel metal1 182 -48 182 -48 1 gnd
rlabel metal1 182 26 182 26 5 vdd
rlabel metal1 172 -6 172 -6 3 A
rlabel metal1 193 -6 193 -6 7 Z
<< end >>
