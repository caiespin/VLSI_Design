magic
tech scmos
timestamp 1552750044
<< nwell >>
rect -4 48 31 105
<< ntransistor >>
rect 7 6 9 33
rect 12 6 14 33
<< ptransistor >>
rect 12 74 14 81
<< ndiffusion >>
rect 6 6 7 33
rect 9 6 12 33
rect 14 6 15 33
<< pdiffusion >>
rect 11 74 12 81
rect 14 74 15 81
<< ndcontact >>
rect 2 6 6 33
rect 15 6 19 33
<< pdcontact >>
rect 7 74 11 81
rect 15 74 19 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 24 -2 28 2
<< nsubstratencontact >>
rect 1 98 5 102
rect 23 98 27 102
<< polysilicon >>
rect 12 81 14 88
rect 12 72 14 74
rect 7 33 9 40
rect 12 33 14 48
rect 7 4 9 6
rect 12 4 14 6
<< polycontact >>
rect 14 84 18 88
rect 8 44 12 48
rect 3 36 7 40
<< metal1 >>
rect -1 102 29 103
rect -1 98 1 102
rect 5 98 23 102
rect 27 98 29 102
rect -1 97 29 98
rect 7 81 11 97
rect 18 84 26 88
rect 15 33 19 74
rect 2 3 6 6
rect 22 3 26 84
rect -1 2 29 3
rect -1 -2 0 2
rect 4 -2 24 2
rect 28 -2 29 2
rect -1 -3 29 -2
<< labels >>
rlabel metal1 8 -1 9 0 1 gnd
rlabel metal1 7 99 8 100 1 vdd
rlabel metal1 17 42 17 42 1 Y
rlabel polycontact 5 38 5 38 1 A
rlabel polycontact 10 46 10 46 1 B
<< end >>
