* NGSPICE file created from ADDER.ext - technology: scmos

.global Vdd Gnd 

.subckt FA COUT gnd CIN vdd
M1000 vdd a_11_n26# COUT vdd pfet w=3.6u l=0.6u
+  ad=29.16p pd=52.2u as=5.4p ps=10.2u
M1001 a_43_2# A a_36_2# vdd pfet w=3.6u l=0.6u
+  ad=6.48p pd=10.8u as=17.28p ps=31.2u
M1002 a_11_n26# B a_43_2# vdd pfet w=3.6u l=0.6u
+  ad=6.48p pd=10.8u as=0p ps=0u
M1003 a_36_2# CIN a_11_n26# vdd pfet w=3.6u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1004 vdd A a_36_2# vdd pfet w=3.6u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_36_2# B vdd vdd pfet w=3.6u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_105_2# A vdd vdd pfet w=3.6u l=0.6u
+  ad=18.36p pd=31.8u as=0p ps=0u
M1007 vdd B a_105_2# vdd pfet w=3.6u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_105_2# CIN vdd vdd pfet w=3.6u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_129_2# A a_105_2# vdd pfet w=3.6u l=0.6u
+  ad=6.48p pd=10.8u as=0p ps=0u
M1010 a_137_2# B a_129_2# vdd pfet w=3.6u l=0.6u
+  ad=6.48p pd=10.8u as=0p ps=0u
M1011 a_98_n43# CIN a_137_2# vdd pfet w=3.6u l=0.6u
+  ad=6.48p pd=10.8u as=0p ps=0u
M1012 a_105_2# a_11_n26# a_98_n43# vdd pfet w=3.6u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1013 SUM a_98_n43# vdd vdd pfet w=3.6u l=0.6u
+  ad=5.4p pd=10.2u as=0p ps=0u
M1014 gnd a_11_n26# COUT Gnd nfet w=1.2u l=0.6u
+  ad=11.88p pd=34.2u as=1.8p ps=5.4u
M1015 SUM a_98_n43# gnd Gnd nfet w=1.2u l=0.6u
+  ad=1.8p pd=5.4u as=0p ps=0u
M1016 gnd A a_36_n43# Gnd nfet w=1.2u l=0.6u
+  ad=0p pd=0u as=3.96p ps=11.4u
M1017 a_36_n43# B gnd Gnd nfet w=1.2u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_11_n26# CIN a_36_n43# Gnd nfet w=1.2u l=0.6u
+  ad=2.16p pd=6u as=0p ps=0u
M1019 a_67_n43# A a_11_n26# Gnd nfet w=1.2u l=0.6u
+  ad=2.16p pd=6u as=0p ps=0u
M1020 gnd B a_67_n43# Gnd nfet w=1.2u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_105_n43# A a_98_n43# Gnd nfet w=1.2u l=0.6u
+  ad=2.16p pd=6u as=3.6p ps=10.8u
M1022 a_113_n43# B a_105_n43# Gnd nfet w=1.2u l=0.6u
+  ad=2.16p pd=6u as=0p ps=0u
M1023 gnd CIN a_113_n43# Gnd nfet w=1.2u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_129_n43# A gnd Gnd nfet w=1.2u l=0.6u
+  ad=4.32p pd=12u as=0p ps=0u
M1025 gnd B a_129_n43# Gnd nfet w=1.2u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_129_n43# CIN gnd Gnd nfet w=1.2u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_98_n43# a_11_n26# a_129_n43# Gnd nfet w=1.2u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
.ends


* Top level circuit ADDER

XFA_7 FA_7/COUT FA_0/gnd FA_7/CIN FA_0/vdd FA
XFA_6 FA_7/CIN FA_0/gnd FA_6/CIN FA_0/vdd FA
XFA_5 FA_6/CIN FA_0/gnd FA_5/CIN FA_0/vdd FA
XFA_4 FA_5/CIN FA_0/gnd FA_4/CIN FA_0/vdd FA
XFA_3 FA_4/CIN FA_0/gnd FA_3/CIN FA_0/vdd FA
XFA_2 FA_3/CIN FA_0/gnd FA_2/CIN FA_0/vdd FA
XFA_1 FA_2/CIN FA_0/gnd FA_1/CIN FA_0/vdd FA
XFA_0 FA_1/CIN FA_0/gnd FA_0/CIN FA_0/vdd FA
.end

