magic
tech scmos
timestamp 1552751125
<< nwell >>
rect -8 53 24 105
<< ntransistor >>
rect 7 6 9 19
rect 15 6 17 19
<< ptransistor >>
rect 7 59 9 66
<< ndiffusion >>
rect 6 6 7 19
rect 9 6 10 19
rect 14 6 15 19
rect 17 6 18 19
<< pdiffusion >>
rect 6 59 7 66
rect 9 59 10 66
<< ndcontact >>
rect 2 6 6 19
rect 10 6 14 19
rect 18 6 22 19
<< pdcontact >>
rect 2 59 6 66
rect 10 59 14 66
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 66 9 68
rect 7 52 9 59
rect 7 19 9 26
rect 15 19 17 33
rect 7 4 9 6
rect 15 4 17 6
<< polycontact >>
rect 3 52 7 56
rect 3 22 7 26
rect 17 29 21 33
<< metal1 >>
rect -7 102 23 103
rect -7 98 -2 102
rect 2 98 14 102
rect 18 98 23 102
rect -7 97 23 98
rect 2 66 6 97
rect -5 52 3 56
rect -5 3 -1 52
rect 10 19 14 59
rect 2 3 6 6
rect 18 3 22 6
rect -7 2 23 3
rect -7 -2 -2 2
rect 2 -2 14 2
rect 18 -2 23 2
rect -7 -3 23 -2
<< labels >>
rlabel metal1 9 0 9 0 1 GND
rlabel metal1 11 100 11 100 5 VDD
rlabel metal1 12 38 12 38 1 Y
rlabel polycontact 5 24 5 24 1 A
rlabel polycontact 19 31 19 31 7 B
<< end >>
