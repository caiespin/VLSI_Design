* SPICE3 file created from NOR2X1_new.ext - technology: scmos

.subckt NOR2X1_new A B Y vdd gnd
M1000 Y GND VDD VDD pfet w=2.1u l=0.6u
+  ad=3.15p pd=7.2u as=3.15p ps=7.2u
M1001 Y A GND Gnd nfet w=3.9u l=0.6u
+  ad=7.02p pd=11.4u as=11.7p ps=21.6u
M1002 GND B Y Gnd nfet w=3.9u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
C0 GND Gnd 5.83fF
C1 VDD Gnd 5.84fF
.ends

X100 A B Z VDD GND NOR2X1_new
.end