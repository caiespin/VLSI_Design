magic
tech scmos
timestamp 1550209003
<< metal1 >>
rect -79 73 1515 77
rect 161 33 173 36
rect 361 33 373 36
rect 561 33 573 36
rect 761 33 773 36
rect 961 33 973 36
rect 1161 33 1173 36
rect 1361 33 1369 36
rect -79 0 1515 4
<< m2contact >>
rect 105 32 109 36
rect 157 32 161 36
rect 305 32 309 36
rect 357 32 361 36
rect 505 32 509 36
rect 557 32 561 36
rect 705 32 709 36
rect 757 32 761 36
rect 905 32 909 36
rect 957 32 961 36
rect 1105 32 1109 36
rect 1157 32 1161 36
rect 1305 32 1309 36
rect 1357 32 1361 36
<< metal2 >>
rect 109 32 157 36
rect 309 32 357 36
rect 509 32 557 36
rect 709 32 757 36
rect 909 32 957 36
rect 1109 32 1157 36
rect 1309 32 1357 36
use FA  FA_0
timestamp 1550166721
transform -1 0 115 0 1 50
box 0 -50 194 27
use FA  FA_1
timestamp 1550166721
transform -1 0 315 0 1 50
box 0 -50 194 27
use FA  FA_2
timestamp 1550166721
transform -1 0 515 0 1 50
box 0 -50 194 27
use FA  FA_3
timestamp 1550166721
transform -1 0 715 0 1 50
box 0 -50 194 27
use FA  FA_4
timestamp 1550166721
transform -1 0 915 0 1 50
box 0 -50 194 27
use FA  FA_5
timestamp 1550166721
transform -1 0 1115 0 1 50
box 0 -50 194 27
use FA  FA_6
timestamp 1550166721
transform -1 0 1315 0 1 50
box 0 -50 194 27
use FA  FA_7
timestamp 1550166721
transform -1 0 1515 0 1 50
box 0 -50 194 27
<< end >>
